library verilog;
use verilog.vl_types.all;
entity view_vlg_vec_tst is
end view_vlg_vec_tst;
