library verilog;
use verilog.vl_types.all;
entity tb_f_word_set is
end tb_f_word_set;
