library verilog;
use verilog.vl_types.all;
entity tb_dds is
end tb_dds;
